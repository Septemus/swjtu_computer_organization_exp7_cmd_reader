library verilog;
use verilog.vl_types.all;
entity exp7_vlg_vec_tst is
end exp7_vlg_vec_tst;
